-------------------------------------------------------------------------------
--
-- Title       : forwarding_mux
-- Design      : alu
-- Author      : Michael
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : C:/Users/Michael/Desktop/Stony Brook University/Fall 2024/ESE 345/Project/ESE_345_Project/alu/src/forwarding_mux.vhd
-- Generated   : Thu Nov 28 21:30:42 2024
-- From        : Interface description file
-- By          : ItfToHdl ver. 1.0
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--    and may be overwritten
--{entity {forwarding_mux} architecture {behavior}}

library ieee;
use ieee.std_logic_1164.all;

entity forwarding_mux is
	port(
	fwd_reg1, fwd_reg2, fwd_reg3 : in std_logic
	
	);
end forwarding_mux;

--}} End of automatically maintained section

architecture behavior of forwarding_mux is
begin

	-- Enter your statements here --

end behavior;
